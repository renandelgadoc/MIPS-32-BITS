library verilog;
use verilog.vl_types.all;
entity OAC_Lab2_vlg_vec_tst is
end OAC_Lab2_vlg_vec_tst;
